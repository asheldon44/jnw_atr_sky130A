magic
tech sky130A
magscale 1 1
timestamp 1723932000
<< checkpaint >>
rect 0 0 576 400
<< pdiff >>
rect 208 20 368 60
rect 208 60 368 100
rect 208 100 368 140
rect 208 140 368 180
rect 208 180 368 220
rect 208 220 368 260
rect 208 260 368 300
rect 208 300 368 340
rect 208 340 368 380
<< ntap >>
rect -48 -20 48 20
rect 528 -20 624 20
rect -48 20 48 60
rect 528 20 624 60
rect -48 60 48 100
rect 528 60 624 100
rect -48 100 48 140
rect 528 100 624 140
rect -48 140 48 180
rect 528 140 624 180
rect -48 180 48 220
rect 528 180 624 220
rect -48 220 48 260
rect 528 220 624 260
rect -48 260 48 300
rect 528 260 624 300
rect -48 300 48 340
rect 528 300 624 340
rect -48 340 48 380
rect 528 340 624 380
rect -48 380 48 420
rect 528 380 624 420
<< poly >>
rect 80 73 496 167
rect 80 233 496 327
rect 80 -11 496 11
rect 80 100 112 140
rect 464 100 496 140
rect 80 140 112 180
rect 464 140 496 180
rect 80 180 112 220
rect 464 180 496 220
rect 80 220 112 260
rect 464 220 496 260
rect 80 260 112 300
rect 464 260 496 300
rect 80 389 496 411
<< m1 >>
rect 80 180 112 220
rect 144 300 240 340
rect 336 20 432 60
rect 80 20 112 60
rect 144 20 240 60
rect 336 20 432 60
rect 80 60 112 100
rect 144 60 240 100
rect 336 60 432 100
rect 80 100 112 140
rect 144 100 240 140
rect 336 100 432 140
rect 80 140 112 180
rect 144 140 240 180
rect 336 140 432 180
rect 80 180 112 220
rect 144 180 240 220
rect 336 180 432 220
rect 80 220 112 260
rect 144 220 240 260
rect 336 220 432 260
rect 80 260 112 300
rect 144 260 240 300
rect 336 260 432 300
rect 80 300 112 340
rect 144 300 240 340
rect 336 300 432 340
rect 80 340 112 380
rect 144 340 240 380
rect 336 340 432 380
<< pcontact >>
rect 85 150 106 160
rect 85 160 106 170
rect 85 170 106 180
rect 469 150 490 160
rect 469 160 490 170
rect 469 170 490 180
rect 85 180 106 190
rect 85 190 106 200
rect 85 200 106 210
rect 85 210 106 220
rect 469 180 490 190
rect 469 190 490 200
rect 469 200 490 210
rect 469 210 490 220
rect 85 220 106 230
rect 85 230 106 240
rect 85 240 106 250
rect 469 220 490 230
rect 469 230 490 240
rect 469 240 490 250
<< locali >>
rect -48 -20 48 20
rect 528 -20 624 20
rect -48 20 48 60
rect 144 20 368 60
rect 528 20 624 60
rect -48 60 48 100
rect 528 60 624 100
rect -48 100 48 140
rect 528 100 624 140
rect -48 140 48 180
rect 80 140 112 180
rect 464 140 496 180
rect 528 140 624 180
rect -48 180 48 220
rect -48 180 48 220
rect 80 180 112 220
rect 208 180 432 220
rect 464 180 496 220
rect 528 180 624 220
rect -48 220 48 260
rect 80 220 112 260
rect 464 220 496 260
rect 528 220 624 260
rect -48 260 48 300
rect 528 260 624 300
rect -48 300 48 340
rect 528 300 624 340
rect -48 340 48 380
rect 144 340 368 380
rect 528 340 624 380
rect -48 380 48 420
rect 528 380 624 420
<< ntapc >>
rect -16 100 16 140
rect 560 100 592 140
rect -16 140 16 180
rect 560 140 592 180
rect -16 180 16 220
rect 560 180 592 220
rect -16 220 16 260
rect 560 220 592 260
rect -16 260 16 300
rect 560 260 592 300
<< pdcontact >>
rect 224 30 240 40
rect 224 40 240 50
rect 240 30 272 40
rect 240 40 272 50
rect 272 30 304 40
rect 272 40 304 50
rect 304 30 336 40
rect 304 40 336 50
rect 336 30 352 40
rect 336 40 352 50
rect 224 190 240 200
rect 224 200 240 210
rect 240 190 272 200
rect 240 200 272 210
rect 272 190 304 200
rect 272 200 304 210
rect 304 190 336 200
rect 304 200 336 210
rect 336 190 352 200
rect 336 200 352 210
rect 224 350 240 360
rect 224 360 240 370
rect 240 350 272 360
rect 240 360 272 370
rect 272 350 304 360
rect 272 360 304 370
rect 304 350 336 360
rect 304 360 336 370
rect 336 350 352 360
rect 336 360 352 370
<< viali >>
rect 160 24 176 28
rect 160 28 176 32
rect 160 32 176 36
rect 160 36 176 40
rect 160 40 176 44
rect 160 44 176 48
rect 160 48 176 52
rect 160 52 176 56
rect 176 24 208 28
rect 176 28 208 32
rect 176 32 208 36
rect 176 36 208 40
rect 176 40 208 44
rect 176 44 208 48
rect 176 48 208 52
rect 176 52 208 56
rect 208 24 224 28
rect 208 28 224 32
rect 208 32 224 36
rect 208 36 224 40
rect 208 40 224 44
rect 208 44 224 48
rect 208 48 224 52
rect 208 52 224 56
rect 85 150 106 160
rect 85 160 106 170
rect 85 170 106 180
rect 85 180 106 190
rect 85 190 106 200
rect 85 200 106 210
rect 85 210 106 220
rect 352 184 368 188
rect 352 188 368 192
rect 352 192 368 196
rect 352 196 368 200
rect 352 200 368 204
rect 352 204 368 208
rect 352 208 368 212
rect 352 212 368 216
rect 368 184 400 188
rect 368 188 400 192
rect 368 192 400 196
rect 368 196 400 200
rect 368 200 400 204
rect 368 204 400 208
rect 368 208 400 212
rect 368 212 400 216
rect 400 184 416 188
rect 400 188 416 192
rect 400 192 416 196
rect 400 196 416 200
rect 400 200 416 204
rect 400 204 416 208
rect 400 208 416 212
rect 400 212 416 216
rect 85 220 106 230
rect 85 230 106 240
rect 85 240 106 250
rect 160 344 176 348
rect 160 348 176 352
rect 160 352 176 356
rect 160 356 176 360
rect 160 360 176 364
rect 160 364 176 368
rect 160 368 176 372
rect 160 372 176 376
rect 176 344 208 348
rect 176 348 208 352
rect 176 352 208 356
rect 176 356 208 360
rect 176 360 208 364
rect 176 364 208 368
rect 176 368 208 372
rect 176 372 208 376
rect 208 344 224 348
rect 208 348 224 352
rect 208 352 224 356
rect 208 356 224 360
rect 208 360 224 364
rect 208 364 224 368
rect 208 368 224 372
rect 208 372 224 376
<< nwell >>
rect -92 -64 668 464
<< labels >>
flabel m1 s 80 180 112 220 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel m1 s 144 300 240 340 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s -48 180 48 220 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel m1 s 336 20 432 60 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 576 400
<< end >>
