magic
tech sky130A
magscale 1 1
timestamp 1723932000
<< checkpaint >>
rect 0 0 832 400
<< pdiff >>
rect 208 100 624 140
rect 208 140 624 180
rect 208 180 624 220
rect 208 220 624 260
rect 208 260 624 300
<< ntap >>
rect -48 -20 48 20
rect 784 -20 880 20
rect -48 20 48 60
rect 784 20 880 60
rect -48 60 48 100
rect 784 60 880 100
rect -48 100 48 140
rect 784 100 880 140
rect -48 140 48 180
rect 784 140 880 180
rect -48 180 48 220
rect 784 180 880 220
rect -48 220 48 260
rect 784 220 880 260
rect -48 260 48 300
rect 784 260 880 300
rect -48 300 48 340
rect 784 300 880 340
rect -48 340 48 380
rect 784 340 880 380
rect -48 380 48 420
rect 784 380 880 420
<< poly >>
rect 80 -11 752 11
rect 80 69 752 91
rect 80 149 752 171
rect 80 229 752 251
rect 80 309 752 331
rect 80 389 752 411
rect 80 140 112 180
rect 720 140 752 180
rect 80 180 112 220
rect 720 180 752 220
rect 80 220 112 260
rect 720 220 752 260
<< m1 >>
rect 80 180 112 220
rect 144 300 240 340
rect 592 20 688 60
rect 80 20 112 60
rect 144 20 240 60
rect 592 20 688 60
rect 80 60 112 100
rect 144 60 240 100
rect 592 60 688 100
rect 80 100 112 140
rect 144 100 240 140
rect 592 100 688 140
rect 80 140 112 180
rect 144 140 240 180
rect 592 140 688 180
rect 80 180 112 220
rect 144 180 240 220
rect 592 180 688 220
rect 80 220 112 260
rect 144 220 240 260
rect 592 220 688 260
rect 80 260 112 300
rect 144 260 240 300
rect 592 260 688 300
rect 80 300 112 340
rect 144 300 240 340
rect 592 300 688 340
rect 80 340 112 380
rect 144 340 240 380
rect 592 340 688 380
<< pcontact >>
rect 85 150 106 160
rect 85 160 106 170
rect 85 170 106 180
rect 725 150 746 160
rect 725 160 746 170
rect 725 170 746 180
rect 85 180 106 190
rect 85 190 106 200
rect 85 200 106 210
rect 85 210 106 220
rect 725 180 746 190
rect 725 190 746 200
rect 725 200 746 210
rect 725 210 746 220
rect 85 220 106 230
rect 85 230 106 240
rect 85 240 106 250
rect 725 220 746 230
rect 725 230 746 240
rect 725 240 746 250
<< locali >>
rect -48 -20 48 20
rect 784 -20 880 20
rect -48 20 48 60
rect 784 20 880 60
rect -48 60 48 100
rect 784 60 880 100
rect -48 100 48 140
rect 144 100 624 140
rect 784 100 880 140
rect -48 140 48 180
rect 80 140 112 180
rect 720 140 752 180
rect 784 140 880 180
rect -48 180 48 220
rect -48 180 48 220
rect 80 180 112 220
rect 208 180 688 220
rect 720 180 752 220
rect 784 180 880 220
rect -48 220 48 260
rect 80 220 112 260
rect 720 220 752 260
rect 784 220 880 260
rect -48 260 48 300
rect 144 260 624 300
rect 784 260 880 300
rect -48 300 48 340
rect 784 300 880 340
rect -48 340 48 380
rect 784 340 880 380
rect -48 380 48 420
rect 784 380 880 420
<< ntapc >>
rect -16 100 16 140
rect 816 100 848 140
rect -16 140 16 180
rect 816 140 848 180
rect -16 180 16 220
rect 816 180 848 220
rect -16 220 16 260
rect 816 220 848 260
rect -16 260 16 300
rect 816 260 848 300
<< pdcontact >>
rect 224 110 240 120
rect 224 120 240 130
rect 240 110 272 120
rect 240 120 272 130
rect 272 110 304 120
rect 272 120 304 130
rect 304 110 336 120
rect 304 120 336 130
rect 336 110 368 120
rect 336 120 368 130
rect 368 110 400 120
rect 368 120 400 130
rect 400 110 432 120
rect 400 120 432 130
rect 432 110 464 120
rect 432 120 464 130
rect 464 110 496 120
rect 464 120 496 130
rect 496 110 528 120
rect 496 120 528 130
rect 528 110 560 120
rect 528 120 560 130
rect 560 110 592 120
rect 560 120 592 130
rect 592 110 608 120
rect 592 120 608 130
rect 224 190 240 200
rect 224 200 240 210
rect 240 190 272 200
rect 240 200 272 210
rect 272 190 304 200
rect 272 200 304 210
rect 304 190 336 200
rect 304 200 336 210
rect 336 190 368 200
rect 336 200 368 210
rect 368 190 400 200
rect 368 200 400 210
rect 400 190 432 200
rect 400 200 432 210
rect 432 190 464 200
rect 432 200 464 210
rect 464 190 496 200
rect 464 200 496 210
rect 496 190 528 200
rect 496 200 528 210
rect 528 190 560 200
rect 528 200 560 210
rect 560 190 592 200
rect 560 200 592 210
rect 592 190 608 200
rect 592 200 608 210
rect 224 270 240 280
rect 224 280 240 290
rect 240 270 272 280
rect 240 280 272 290
rect 272 270 304 280
rect 272 280 304 290
rect 304 270 336 280
rect 304 280 336 290
rect 336 270 368 280
rect 336 280 368 290
rect 368 270 400 280
rect 368 280 400 290
rect 400 270 432 280
rect 400 280 432 290
rect 432 270 464 280
rect 432 280 464 290
rect 464 270 496 280
rect 464 280 496 290
rect 496 270 528 280
rect 496 280 528 290
rect 528 270 560 280
rect 528 280 560 290
rect 560 270 592 280
rect 560 280 592 290
rect 592 270 608 280
rect 592 280 608 290
<< viali >>
rect 160 104 176 108
rect 160 108 176 112
rect 160 112 176 116
rect 160 116 176 120
rect 160 120 176 124
rect 160 124 176 128
rect 160 128 176 132
rect 160 132 176 136
rect 176 104 208 108
rect 176 108 208 112
rect 176 112 208 116
rect 176 116 208 120
rect 176 120 208 124
rect 176 124 208 128
rect 176 128 208 132
rect 176 132 208 136
rect 208 104 224 108
rect 208 108 224 112
rect 208 112 224 116
rect 208 116 224 120
rect 208 120 224 124
rect 208 124 224 128
rect 208 128 224 132
rect 208 132 224 136
rect 85 150 106 160
rect 85 160 106 170
rect 85 170 106 180
rect 85 180 106 190
rect 85 190 106 200
rect 85 200 106 210
rect 85 210 106 220
rect 608 184 624 188
rect 608 188 624 192
rect 608 192 624 196
rect 608 196 624 200
rect 608 200 624 204
rect 608 204 624 208
rect 608 208 624 212
rect 608 212 624 216
rect 624 184 656 188
rect 624 188 656 192
rect 624 192 656 196
rect 624 196 656 200
rect 624 200 656 204
rect 624 204 656 208
rect 624 208 656 212
rect 624 212 656 216
rect 656 184 672 188
rect 656 188 672 192
rect 656 192 672 196
rect 656 196 672 200
rect 656 200 672 204
rect 656 204 672 208
rect 656 208 672 212
rect 656 212 672 216
rect 85 220 106 230
rect 85 230 106 240
rect 85 240 106 250
rect 160 264 176 268
rect 160 268 176 272
rect 160 272 176 276
rect 160 276 176 280
rect 160 280 176 284
rect 160 284 176 288
rect 160 288 176 292
rect 160 292 176 296
rect 176 264 208 268
rect 176 268 208 272
rect 176 272 208 276
rect 176 276 208 280
rect 176 280 208 284
rect 176 284 208 288
rect 176 288 208 292
rect 176 292 208 296
rect 208 264 224 268
rect 208 268 224 272
rect 208 272 224 276
rect 208 276 224 280
rect 208 280 224 284
rect 208 284 224 288
rect 208 288 224 292
rect 208 292 224 296
<< nwell >>
rect -92 -64 924 464
<< labels >>
flabel m1 s 80 180 112 220 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel m1 s 144 300 240 340 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s -48 180 48 220 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel m1 s 592 20 688 60 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 832 400
<< end >>
