
//-------------------------------------------------------------
// JNWATR_PCH_2C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module JNWATR_PCH_2C1F2(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// JNWATR_PCH_2C5F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module JNWATR_PCH_2C5F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// JNWATR_PCH_4C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module JNWATR_PCH_4C1F2(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// JNWATR_PCH_4C5F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module JNWATR_PCH_4C5F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// JNWATR_PCH_8C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module JNWATR_PCH_8C1F2(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// JNWATR_PCH_8C5F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module JNWATR_PCH_8C5F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// JNWATR_PCH_12C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module JNWATR_PCH_12C1F2(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// JNWATR_PCH_12C5F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module JNWATR_PCH_12C5F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// JNWATR_NCH_2C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module JNWATR_NCH_2C1F2(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// JNWATR_NCH_2C5F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module JNWATR_NCH_2C5F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// JNWATR_NCH_4C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module JNWATR_NCH_4C1F2(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// JNWATR_NCH_4C5F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module JNWATR_NCH_4C5F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// JNWATR_NCH_8C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module JNWATR_NCH_8C1F2(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// JNWATR_NCH_8C5F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module JNWATR_NCH_8C5F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// JNWATR_NCH_12C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module JNWATR_NCH_12C1F2(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// JNWATR_NCH_12C5F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module JNWATR_NCH_12C5F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule
