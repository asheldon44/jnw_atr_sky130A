magic
tech sky130B
magscale 1 1
timestamp 1712527200
<< checkpaint >>
rect 0 0 576 400
<< pdiff >>
rect 208 100 368 140
rect 208 140 368 180
rect 208 180 368 220
rect 208 220 368 260
rect 208 260 368 300
<< ntap >>
rect -48 -20 48 20
rect 528 -20 624 20
rect -48 20 48 60
rect 528 20 624 60
rect -48 60 48 100
rect 528 60 624 100
rect -48 100 48 140
rect 528 100 624 140
rect -48 140 48 180
rect 528 140 624 180
rect -48 180 48 220
rect 528 180 624 220
rect -48 220 48 260
rect 528 220 624 260
rect -48 260 48 300
rect 528 260 624 300
rect -48 300 48 340
rect 528 300 624 340
rect -48 340 48 380
rect 528 340 624 380
rect -48 380 48 420
rect 528 380 624 420
<< poly >>
rect 80 -11 496 11
rect 80 69 496 91
rect 80 149 496 171
rect 80 229 496 251
rect 80 309 496 331
rect 80 389 496 411
rect 80 140 112 180
rect 464 140 496 180
rect 80 180 112 220
rect 464 180 496 220
rect 80 220 112 260
rect 464 220 496 260
<< m1 >>
rect 80 180 112 220
rect 144 300 240 340
rect 336 20 432 60
rect 80 20 112 60
rect 144 20 240 60
rect 336 20 432 60
rect 80 60 112 100
rect 144 60 240 100
rect 336 60 432 100
rect 80 100 112 140
rect 144 100 240 140
rect 336 100 432 140
rect 80 140 112 180
rect 144 140 240 180
rect 336 140 432 180
rect 80 180 112 220
rect 144 180 240 220
rect 336 180 432 220
rect 80 220 112 260
rect 144 220 240 260
rect 336 220 432 260
rect 80 260 112 300
rect 144 260 240 300
rect 336 260 432 300
rect 80 300 112 340
rect 144 300 240 340
rect 336 300 432 340
rect 80 340 112 380
rect 144 340 240 380
rect 336 340 432 380
<< pcontact >>
rect 85 150 106 160
rect 85 160 106 170
rect 85 170 106 180
rect 469 150 490 160
rect 469 160 490 170
rect 469 170 490 180
rect 85 180 106 190
rect 85 190 106 200
rect 85 200 106 210
rect 85 210 106 220
rect 469 180 490 190
rect 469 190 490 200
rect 469 200 490 210
rect 469 210 490 220
rect 85 220 106 230
rect 85 230 106 240
rect 85 240 106 250
rect 469 220 490 230
rect 469 230 490 240
rect 469 240 490 250
<< locali >>
rect -48 -20 48 20
rect 528 -20 624 20
rect -48 20 48 60
rect 528 20 624 60
rect -48 60 48 100
rect 528 60 624 100
rect -48 100 48 140
rect 144 100 368 140
rect 528 100 624 140
rect -48 140 48 180
rect 80 140 112 180
rect 464 140 496 180
rect 528 140 624 180
rect -48 180 48 220
rect -48 180 48 220
rect 80 180 112 220
rect 208 180 432 220
rect 464 180 496 220
rect 528 180 624 220
rect -48 220 48 260
rect 80 220 112 260
rect 464 220 496 260
rect 528 220 624 260
rect -48 260 48 300
rect 144 260 368 300
rect 528 260 624 300
rect -48 300 48 340
rect 528 300 624 340
rect -48 340 48 380
rect 528 340 624 380
rect -48 380 48 420
rect 528 380 624 420
<< ntapc >>
rect -16 100 16 140
rect 560 100 592 140
rect -16 140 16 180
rect 560 140 592 180
rect -16 180 16 220
rect 560 180 592 220
rect -16 220 16 260
rect 560 220 592 260
rect -16 260 16 300
rect 560 260 592 300
<< pdcontact >>
rect 224 110 240 120
rect 224 120 240 130
rect 240 110 272 120
rect 240 120 272 130
rect 272 110 304 120
rect 272 120 304 130
rect 304 110 336 120
rect 304 120 336 130
rect 336 110 352 120
rect 336 120 352 130
rect 224 190 240 200
rect 224 200 240 210
rect 240 190 272 200
rect 240 200 272 210
rect 272 190 304 200
rect 272 200 304 210
rect 304 190 336 200
rect 304 200 336 210
rect 336 190 352 200
rect 336 200 352 210
rect 224 270 240 280
rect 224 280 240 290
rect 240 270 272 280
rect 240 280 272 290
rect 272 270 304 280
rect 272 280 304 290
rect 304 270 336 280
rect 304 280 336 290
rect 336 270 352 280
rect 336 280 352 290
<< viali >>
rect 160 104 176 108
rect 160 108 176 112
rect 160 112 176 116
rect 160 116 176 120
rect 160 120 176 124
rect 160 124 176 128
rect 160 128 176 132
rect 160 132 176 136
rect 176 104 208 108
rect 176 108 208 112
rect 176 112 208 116
rect 176 116 208 120
rect 176 120 208 124
rect 176 124 208 128
rect 176 128 208 132
rect 176 132 208 136
rect 208 104 224 108
rect 208 108 224 112
rect 208 112 224 116
rect 208 116 224 120
rect 208 120 224 124
rect 208 124 224 128
rect 208 128 224 132
rect 208 132 224 136
rect 85 150 106 160
rect 85 160 106 170
rect 85 170 106 180
rect 85 180 106 190
rect 85 190 106 200
rect 85 200 106 210
rect 85 210 106 220
rect 352 184 368 188
rect 352 188 368 192
rect 352 192 368 196
rect 352 196 368 200
rect 352 200 368 204
rect 352 204 368 208
rect 352 208 368 212
rect 352 212 368 216
rect 368 184 400 188
rect 368 188 400 192
rect 368 192 400 196
rect 368 196 400 200
rect 368 200 400 204
rect 368 204 400 208
rect 368 208 400 212
rect 368 212 400 216
rect 400 184 416 188
rect 400 188 416 192
rect 400 192 416 196
rect 400 196 416 200
rect 400 200 416 204
rect 400 204 416 208
rect 400 208 416 212
rect 400 212 416 216
rect 85 220 106 230
rect 85 230 106 240
rect 85 240 106 250
rect 160 264 176 268
rect 160 268 176 272
rect 160 272 176 276
rect 160 276 176 280
rect 160 280 176 284
rect 160 284 176 288
rect 160 288 176 292
rect 160 292 176 296
rect 176 264 208 268
rect 176 268 208 272
rect 176 272 208 276
rect 176 276 208 280
rect 176 280 208 284
rect 176 284 208 288
rect 176 288 208 292
rect 176 292 208 296
rect 208 264 224 268
rect 208 268 224 272
rect 208 272 224 276
rect 208 276 224 280
rect 208 280 224 284
rect 208 284 224 288
rect 208 288 224 292
rect 208 292 224 296
<< nwell >>
rect -92 -64 668 464
<< labels >>
flabel m1 s 80 180 112 220 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel m1 s 144 300 240 340 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s -48 180 48 220 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel m1 s 336 20 432 60 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 576 400
<< end >>
