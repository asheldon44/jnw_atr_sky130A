magic
tech sky130A
magscale 1 1
timestamp 1723932000
<< checkpaint >>
rect 0 0 512 400
<< pdiff >>
rect 208 100 304 140
rect 208 140 304 180
rect 208 180 304 220
rect 208 220 304 260
rect 208 260 304 300
<< ntap >>
rect -48 -20 48 20
rect 464 -20 560 20
rect -48 20 48 60
rect 464 20 560 60
rect -48 60 48 100
rect 464 60 560 100
rect -48 100 48 140
rect 464 100 560 140
rect -48 140 48 180
rect 464 140 560 180
rect -48 180 48 220
rect 464 180 560 220
rect -48 220 48 260
rect 464 220 560 260
rect -48 260 48 300
rect 464 260 560 300
rect -48 300 48 340
rect 464 300 560 340
rect -48 340 48 380
rect 464 340 560 380
rect -48 380 48 420
rect 464 380 560 420
<< poly >>
rect 80 -11 432 11
rect 80 69 432 91
rect 80 149 432 171
rect 80 229 432 251
rect 80 309 432 331
rect 80 389 432 411
rect 80 140 112 180
rect 400 140 432 180
rect 80 180 112 220
rect 400 180 432 220
rect 80 220 112 260
rect 400 220 432 260
<< m1 >>
rect 80 180 112 220
rect 144 300 240 340
rect 272 20 368 60
rect 80 20 112 60
rect 144 20 240 60
rect 272 20 368 60
rect 80 60 112 100
rect 144 60 240 100
rect 272 60 368 100
rect 80 100 112 140
rect 144 100 240 140
rect 272 100 368 140
rect 80 140 112 180
rect 144 140 240 180
rect 272 140 368 180
rect 80 180 112 220
rect 144 180 240 220
rect 272 180 368 220
rect 80 220 112 260
rect 144 220 240 260
rect 272 220 368 260
rect 80 260 112 300
rect 144 260 240 300
rect 272 260 368 300
rect 80 300 112 340
rect 144 300 240 340
rect 272 300 368 340
rect 80 340 112 380
rect 144 340 240 380
rect 272 340 368 380
<< pcontact >>
rect 85 150 106 160
rect 85 160 106 170
rect 85 170 106 180
rect 405 150 426 160
rect 405 160 426 170
rect 405 170 426 180
rect 85 180 106 190
rect 85 190 106 200
rect 85 200 106 210
rect 85 210 106 220
rect 405 180 426 190
rect 405 190 426 200
rect 405 200 426 210
rect 405 210 426 220
rect 85 220 106 230
rect 85 230 106 240
rect 85 240 106 250
rect 405 220 426 230
rect 405 230 426 240
rect 405 240 426 250
<< locali >>
rect -48 -20 48 20
rect 464 -20 560 20
rect -48 20 48 60
rect 464 20 560 60
rect -48 60 48 100
rect 464 60 560 100
rect -48 100 48 140
rect 144 100 304 140
rect 464 100 560 140
rect -48 140 48 180
rect 80 140 112 180
rect 400 140 432 180
rect 464 140 560 180
rect -48 180 48 220
rect -48 180 48 220
rect 80 180 112 220
rect 208 180 368 220
rect 400 180 432 220
rect 464 180 560 220
rect -48 220 48 260
rect 80 220 112 260
rect 400 220 432 260
rect 464 220 560 260
rect -48 260 48 300
rect 144 260 304 300
rect 464 260 560 300
rect -48 300 48 340
rect 464 300 560 340
rect -48 340 48 380
rect 464 340 560 380
rect -48 380 48 420
rect 464 380 560 420
<< ntapc >>
rect -16 100 16 140
rect 496 100 528 140
rect -16 140 16 180
rect 496 140 528 180
rect -16 180 16 220
rect 496 180 528 220
rect -16 220 16 260
rect 496 220 528 260
rect -16 260 16 300
rect 496 260 528 300
<< pdcontact >>
rect 224 110 240 120
rect 224 120 240 130
rect 240 110 272 120
rect 240 120 272 130
rect 272 110 288 120
rect 272 120 288 130
rect 224 190 240 200
rect 224 200 240 210
rect 240 190 272 200
rect 240 200 272 210
rect 272 190 288 200
rect 272 200 288 210
rect 224 270 240 280
rect 224 280 240 290
rect 240 270 272 280
rect 240 280 272 290
rect 272 270 288 280
rect 272 280 288 290
<< viali >>
rect 160 104 176 108
rect 160 108 176 112
rect 160 112 176 116
rect 160 116 176 120
rect 160 120 176 124
rect 160 124 176 128
rect 160 128 176 132
rect 160 132 176 136
rect 176 104 208 108
rect 176 108 208 112
rect 176 112 208 116
rect 176 116 208 120
rect 176 120 208 124
rect 176 124 208 128
rect 176 128 208 132
rect 176 132 208 136
rect 208 104 224 108
rect 208 108 224 112
rect 208 112 224 116
rect 208 116 224 120
rect 208 120 224 124
rect 208 124 224 128
rect 208 128 224 132
rect 208 132 224 136
rect 85 150 106 160
rect 85 160 106 170
rect 85 170 106 180
rect 85 180 106 190
rect 85 190 106 200
rect 85 200 106 210
rect 85 210 106 220
rect 288 184 304 188
rect 288 188 304 192
rect 288 192 304 196
rect 288 196 304 200
rect 288 200 304 204
rect 288 204 304 208
rect 288 208 304 212
rect 288 212 304 216
rect 304 184 336 188
rect 304 188 336 192
rect 304 192 336 196
rect 304 196 336 200
rect 304 200 336 204
rect 304 204 336 208
rect 304 208 336 212
rect 304 212 336 216
rect 336 184 352 188
rect 336 188 352 192
rect 336 192 352 196
rect 336 196 352 200
rect 336 200 352 204
rect 336 204 352 208
rect 336 208 352 212
rect 336 212 352 216
rect 85 220 106 230
rect 85 230 106 240
rect 85 240 106 250
rect 160 264 176 268
rect 160 268 176 272
rect 160 272 176 276
rect 160 276 176 280
rect 160 280 176 284
rect 160 284 176 288
rect 160 288 176 292
rect 160 292 176 296
rect 176 264 208 268
rect 176 268 208 272
rect 176 272 208 276
rect 176 276 208 280
rect 176 280 208 284
rect 176 284 208 288
rect 176 288 208 292
rect 176 292 208 296
rect 208 264 224 268
rect 208 268 224 272
rect 208 272 224 276
rect 208 276 224 280
rect 208 280 224 284
rect 208 284 224 288
rect 208 288 224 292
rect 208 292 224 296
<< nwell >>
rect -92 -64 604 464
<< labels >>
flabel m1 s 80 180 112 220 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel m1 s 144 300 240 340 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s -48 180 48 220 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel m1 s 272 20 368 60 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 512 400
<< end >>
