magic
tech sky130B
magscale 1 1
timestamp 1712527200
<< checkpaint >>
rect 0 0 512 400
<< pdiff >>
rect 208 20 304 60
rect 208 60 304 100
rect 208 100 304 140
rect 208 140 304 180
rect 208 180 304 220
rect 208 220 304 260
rect 208 260 304 300
rect 208 300 304 340
rect 208 340 304 380
<< ptap >>
rect -48 -20 48 20
rect 464 -20 560 20
rect -48 20 48 60
rect 464 20 560 60
rect -48 60 48 100
rect 464 60 560 100
rect -48 100 48 140
rect 464 100 560 140
rect -48 140 48 180
rect 464 140 560 180
rect -48 180 48 220
rect 464 180 560 220
rect -48 220 48 260
rect 464 220 560 260
rect -48 260 48 300
rect 464 260 560 300
rect -48 300 48 340
rect 464 300 560 340
rect -48 340 48 380
rect 464 340 560 380
rect -48 380 48 420
rect 464 380 560 420
<< poly >>
rect 80 73 432 167
rect 80 233 432 327
rect 80 -11 432 11
rect 80 100 112 140
rect 400 100 432 140
rect 80 140 112 180
rect 400 140 432 180
rect 80 180 112 220
rect 400 180 432 220
rect 80 220 112 260
rect 400 220 432 260
rect 80 260 112 300
rect 400 260 432 300
rect 80 389 432 411
<< m1 >>
rect 80 180 112 220
rect 144 300 240 340
rect 272 20 368 60
rect 80 20 112 60
rect 144 20 240 60
rect 272 20 368 60
rect 80 60 112 100
rect 144 60 240 100
rect 272 60 368 100
rect 80 100 112 140
rect 144 100 240 140
rect 272 100 368 140
rect 80 140 112 180
rect 144 140 240 180
rect 272 140 368 180
rect 80 180 112 220
rect 144 180 240 220
rect 272 180 368 220
rect 80 220 112 260
rect 144 220 240 260
rect 272 220 368 260
rect 80 260 112 300
rect 144 260 240 300
rect 272 260 368 300
rect 80 300 112 340
rect 144 300 240 340
rect 272 300 368 340
rect 80 340 112 380
rect 144 340 240 380
rect 272 340 368 380
<< pcontact >>
rect 85 150 106 160
rect 85 160 106 170
rect 85 170 106 180
rect 405 150 426 160
rect 405 160 426 170
rect 405 170 426 180
rect 85 180 106 190
rect 85 190 106 200
rect 85 200 106 210
rect 85 210 106 220
rect 405 180 426 190
rect 405 190 426 200
rect 405 200 426 210
rect 405 210 426 220
rect 85 220 106 230
rect 85 230 106 240
rect 85 240 106 250
rect 405 220 426 230
rect 405 230 426 240
rect 405 240 426 250
<< locali >>
rect -48 -20 48 20
rect 464 -20 560 20
rect -48 20 48 60
rect 144 20 304 60
rect 464 20 560 60
rect -48 60 48 100
rect 464 60 560 100
rect -48 100 48 140
rect 464 100 560 140
rect -48 140 48 180
rect 80 140 112 180
rect 400 140 432 180
rect 464 140 560 180
rect -48 180 48 220
rect -48 180 48 220
rect 80 180 112 220
rect 208 180 368 220
rect 400 180 432 220
rect 464 180 560 220
rect -48 220 48 260
rect 80 220 112 260
rect 400 220 432 260
rect 464 220 560 260
rect -48 260 48 300
rect 464 260 560 300
rect -48 300 48 340
rect 464 300 560 340
rect -48 340 48 380
rect 144 340 304 380
rect 464 340 560 380
rect -48 380 48 420
rect 464 380 560 420
<< ptapc >>
rect -16 100 16 140
rect 496 100 528 140
rect -16 140 16 180
rect 496 140 528 180
rect -16 180 16 220
rect 496 180 528 220
rect -16 220 16 260
rect 496 220 528 260
rect -16 260 16 300
rect 496 260 528 300
<< ndcontact >>
rect 224 30 240 40
rect 224 40 240 50
rect 240 30 272 40
rect 240 40 272 50
rect 272 30 288 40
rect 272 40 288 50
rect 224 190 240 200
rect 224 200 240 210
rect 240 190 272 200
rect 240 200 272 210
rect 272 190 288 200
rect 272 200 288 210
rect 224 350 240 360
rect 224 360 240 370
rect 240 350 272 360
rect 240 360 272 370
rect 272 350 288 360
rect 272 360 288 370
<< viali >>
rect 160 24 176 28
rect 160 28 176 32
rect 160 32 176 36
rect 160 36 176 40
rect 160 40 176 44
rect 160 44 176 48
rect 160 48 176 52
rect 160 52 176 56
rect 176 24 208 28
rect 176 28 208 32
rect 176 32 208 36
rect 176 36 208 40
rect 176 40 208 44
rect 176 44 208 48
rect 176 48 208 52
rect 176 52 208 56
rect 208 24 224 28
rect 208 28 224 32
rect 208 32 224 36
rect 208 36 224 40
rect 208 40 224 44
rect 208 44 224 48
rect 208 48 224 52
rect 208 52 224 56
rect 85 150 106 160
rect 85 160 106 170
rect 85 170 106 180
rect 85 180 106 190
rect 85 190 106 200
rect 85 200 106 210
rect 85 210 106 220
rect 288 184 304 188
rect 288 188 304 192
rect 288 192 304 196
rect 288 196 304 200
rect 288 200 304 204
rect 288 204 304 208
rect 288 208 304 212
rect 288 212 304 216
rect 304 184 336 188
rect 304 188 336 192
rect 304 192 336 196
rect 304 196 336 200
rect 304 200 336 204
rect 304 204 336 208
rect 304 208 336 212
rect 304 212 336 216
rect 336 184 352 188
rect 336 188 352 192
rect 336 192 352 196
rect 336 196 352 200
rect 336 200 352 204
rect 336 204 352 208
rect 336 208 352 212
rect 336 212 352 216
rect 85 220 106 230
rect 85 230 106 240
rect 85 240 106 250
rect 160 344 176 348
rect 160 348 176 352
rect 160 352 176 356
rect 160 356 176 360
rect 160 360 176 364
rect 160 364 176 368
rect 160 368 176 372
rect 160 372 176 376
rect 176 344 208 348
rect 176 348 208 352
rect 176 352 208 356
rect 176 356 208 360
rect 176 360 208 364
rect 176 364 208 368
rect 176 368 208 372
rect 176 372 208 376
rect 208 344 224 348
rect 208 348 224 352
rect 208 352 224 356
rect 208 356 224 360
rect 208 360 224 364
rect 208 364 224 368
rect 208 368 224 372
rect 208 372 224 376
<< pwell >>
rect -92 -64 604 464
<< labels >>
flabel m1 s 80 180 112 220 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel m1 s 144 300 240 340 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s -48 180 48 220 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel m1 s 272 20 368 60 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 512 400
<< end >>
