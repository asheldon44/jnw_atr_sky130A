magic
tech sky130A
magscale 1 1
timestamp 1723932000
<< checkpaint >>
rect 0 0 832 400
<< pdiff >>
rect 208 20 624 60
rect 208 60 624 100
rect 208 100 624 140
rect 208 140 624 180
rect 208 180 624 220
rect 208 220 624 260
rect 208 260 624 300
rect 208 300 624 340
rect 208 340 624 380
<< ptap >>
rect -48 -20 48 20
rect 784 -20 880 20
rect -48 20 48 60
rect 784 20 880 60
rect -48 60 48 100
rect 784 60 880 100
rect -48 100 48 140
rect 784 100 880 140
rect -48 140 48 180
rect 784 140 880 180
rect -48 180 48 220
rect 784 180 880 220
rect -48 220 48 260
rect 784 220 880 260
rect -48 260 48 300
rect 784 260 880 300
rect -48 300 48 340
rect 784 300 880 340
rect -48 340 48 380
rect 784 340 880 380
rect -48 380 48 420
rect 784 380 880 420
<< poly >>
rect 80 73 752 167
rect 80 233 752 327
rect 80 -11 752 11
rect 80 100 112 140
rect 720 100 752 140
rect 80 140 112 180
rect 720 140 752 180
rect 80 180 112 220
rect 720 180 752 220
rect 80 220 112 260
rect 720 220 752 260
rect 80 260 112 300
rect 720 260 752 300
rect 80 389 752 411
<< m1 >>
rect 80 180 112 220
rect 144 300 240 340
rect 592 20 688 60
rect 80 20 112 60
rect 144 20 240 60
rect 592 20 688 60
rect 80 60 112 100
rect 144 60 240 100
rect 592 60 688 100
rect 80 100 112 140
rect 144 100 240 140
rect 592 100 688 140
rect 80 140 112 180
rect 144 140 240 180
rect 592 140 688 180
rect 80 180 112 220
rect 144 180 240 220
rect 592 180 688 220
rect 80 220 112 260
rect 144 220 240 260
rect 592 220 688 260
rect 80 260 112 300
rect 144 260 240 300
rect 592 260 688 300
rect 80 300 112 340
rect 144 300 240 340
rect 592 300 688 340
rect 80 340 112 380
rect 144 340 240 380
rect 592 340 688 380
<< pcontact >>
rect 85 150 106 160
rect 85 160 106 170
rect 85 170 106 180
rect 725 150 746 160
rect 725 160 746 170
rect 725 170 746 180
rect 85 180 106 190
rect 85 190 106 200
rect 85 200 106 210
rect 85 210 106 220
rect 725 180 746 190
rect 725 190 746 200
rect 725 200 746 210
rect 725 210 746 220
rect 85 220 106 230
rect 85 230 106 240
rect 85 240 106 250
rect 725 220 746 230
rect 725 230 746 240
rect 725 240 746 250
<< locali >>
rect -48 -20 48 20
rect 784 -20 880 20
rect -48 20 48 60
rect 144 20 624 60
rect 784 20 880 60
rect -48 60 48 100
rect 784 60 880 100
rect -48 100 48 140
rect 784 100 880 140
rect -48 140 48 180
rect 80 140 112 180
rect 720 140 752 180
rect 784 140 880 180
rect -48 180 48 220
rect -48 180 48 220
rect 80 180 112 220
rect 208 180 688 220
rect 720 180 752 220
rect 784 180 880 220
rect -48 220 48 260
rect 80 220 112 260
rect 720 220 752 260
rect 784 220 880 260
rect -48 260 48 300
rect 784 260 880 300
rect -48 300 48 340
rect 784 300 880 340
rect -48 340 48 380
rect 144 340 624 380
rect 784 340 880 380
rect -48 380 48 420
rect 784 380 880 420
<< ptapc >>
rect -16 100 16 140
rect 816 100 848 140
rect -16 140 16 180
rect 816 140 848 180
rect -16 180 16 220
rect 816 180 848 220
rect -16 220 16 260
rect 816 220 848 260
rect -16 260 16 300
rect 816 260 848 300
<< ndcontact >>
rect 224 30 240 40
rect 224 40 240 50
rect 240 30 272 40
rect 240 40 272 50
rect 272 30 304 40
rect 272 40 304 50
rect 304 30 336 40
rect 304 40 336 50
rect 336 30 368 40
rect 336 40 368 50
rect 368 30 400 40
rect 368 40 400 50
rect 400 30 432 40
rect 400 40 432 50
rect 432 30 464 40
rect 432 40 464 50
rect 464 30 496 40
rect 464 40 496 50
rect 496 30 528 40
rect 496 40 528 50
rect 528 30 560 40
rect 528 40 560 50
rect 560 30 592 40
rect 560 40 592 50
rect 592 30 608 40
rect 592 40 608 50
rect 224 190 240 200
rect 224 200 240 210
rect 240 190 272 200
rect 240 200 272 210
rect 272 190 304 200
rect 272 200 304 210
rect 304 190 336 200
rect 304 200 336 210
rect 336 190 368 200
rect 336 200 368 210
rect 368 190 400 200
rect 368 200 400 210
rect 400 190 432 200
rect 400 200 432 210
rect 432 190 464 200
rect 432 200 464 210
rect 464 190 496 200
rect 464 200 496 210
rect 496 190 528 200
rect 496 200 528 210
rect 528 190 560 200
rect 528 200 560 210
rect 560 190 592 200
rect 560 200 592 210
rect 592 190 608 200
rect 592 200 608 210
rect 224 350 240 360
rect 224 360 240 370
rect 240 350 272 360
rect 240 360 272 370
rect 272 350 304 360
rect 272 360 304 370
rect 304 350 336 360
rect 304 360 336 370
rect 336 350 368 360
rect 336 360 368 370
rect 368 350 400 360
rect 368 360 400 370
rect 400 350 432 360
rect 400 360 432 370
rect 432 350 464 360
rect 432 360 464 370
rect 464 350 496 360
rect 464 360 496 370
rect 496 350 528 360
rect 496 360 528 370
rect 528 350 560 360
rect 528 360 560 370
rect 560 350 592 360
rect 560 360 592 370
rect 592 350 608 360
rect 592 360 608 370
<< viali >>
rect 160 24 176 28
rect 160 28 176 32
rect 160 32 176 36
rect 160 36 176 40
rect 160 40 176 44
rect 160 44 176 48
rect 160 48 176 52
rect 160 52 176 56
rect 176 24 208 28
rect 176 28 208 32
rect 176 32 208 36
rect 176 36 208 40
rect 176 40 208 44
rect 176 44 208 48
rect 176 48 208 52
rect 176 52 208 56
rect 208 24 224 28
rect 208 28 224 32
rect 208 32 224 36
rect 208 36 224 40
rect 208 40 224 44
rect 208 44 224 48
rect 208 48 224 52
rect 208 52 224 56
rect 85 150 106 160
rect 85 160 106 170
rect 85 170 106 180
rect 85 180 106 190
rect 85 190 106 200
rect 85 200 106 210
rect 85 210 106 220
rect 608 184 624 188
rect 608 188 624 192
rect 608 192 624 196
rect 608 196 624 200
rect 608 200 624 204
rect 608 204 624 208
rect 608 208 624 212
rect 608 212 624 216
rect 624 184 656 188
rect 624 188 656 192
rect 624 192 656 196
rect 624 196 656 200
rect 624 200 656 204
rect 624 204 656 208
rect 624 208 656 212
rect 624 212 656 216
rect 656 184 672 188
rect 656 188 672 192
rect 656 192 672 196
rect 656 196 672 200
rect 656 200 672 204
rect 656 204 672 208
rect 656 208 672 212
rect 656 212 672 216
rect 85 220 106 230
rect 85 230 106 240
rect 85 240 106 250
rect 160 344 176 348
rect 160 348 176 352
rect 160 352 176 356
rect 160 356 176 360
rect 160 360 176 364
rect 160 364 176 368
rect 160 368 176 372
rect 160 372 176 376
rect 176 344 208 348
rect 176 348 208 352
rect 176 352 208 356
rect 176 356 208 360
rect 176 360 208 364
rect 176 364 208 368
rect 176 368 208 372
rect 176 372 208 376
rect 208 344 224 348
rect 208 348 224 352
rect 208 352 224 356
rect 208 356 224 360
rect 208 360 224 364
rect 208 364 224 368
rect 208 368 224 372
rect 208 372 224 376
<< pwell >>
rect -92 -64 924 464
<< labels >>
flabel m1 s 80 180 112 220 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel m1 s 144 300 240 340 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s -48 180 48 220 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel m1 s 592 20 688 60 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 832 400
<< end >>
